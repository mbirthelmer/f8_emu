`ifndef F8_OPS_VH_
`define F8_OPS_VH_

`define OP_LR_A_KU		8'h00
`define	OP_LR_A_KL		8'h01
`define OP_LR_A_QU		8'h02
`define OP_LR_A_QL		8'h03
`define OP_LR_KU_A		8'h04
`define OP_LR_KL_A		8'h05
`define OP_LR_QU_A		8'h06
`define OP_LR_QL_A		8'h07
`define OP_LR_K_P		8'h08
`define OP_LR_P_K		8'h09
`define OP_LR_A_IS		8'h0a
`define OP_LR_IS_A		8'h0b
`define OP_PK			8'h0c
`define OP_LR_P0_Q		8'h0d
`define OP_LR_Q_DC		8'h0e
`define OP_LR_DC_Q		8'h0f
`define OP_LR_DC_H		8'h10
`define OP_LR_H_DC		8'h11
`define OP_SR_1			8'h12
`define OP_SL_1			8'h13
`define OP_SR_4			8'h14
`define OP_SL_4			8'h15
`define OP_LM			8'h16
`define OP_ST			8'h17
`define OP_COM			8'h18
`define OP_LNK			8'h19
`define OP_DI			8'h1a
`define OP_EI			8'h1b
`define OP_POP			8'h1c
`define OP_LR_W_J		8'h1d
`define OP_LR_J_W		8'h1e
`define OP_INC			8'h1f
`define OP_LI			8'h20
`define OP_NI			8'h21
`define OP_OI			8'h22
`define OP_XI			8'h23
`define OP_AI			8'h24
`define OP_CI			8'h25
`define OP_IN			8'h26
`define OP_OUT			8'h27
`define OP_PI			8'h28
`define OP_JMP			8'h29
`define OP_DCI			8'h2a
`define OP_NOP			8'h2b
`define OP_XDC			8'h2c
`define OP_DS			8'h3x
`define OP_LR_A_R		8'h4x
`define OP_LR_R_A		8'h5x
`define OP_LISU			8'b01100xxx
`define OP_LISL			8'b01101xxx
`define OP_LIS			8'h7x
`define OP_BT			8'b10000xxx
`define OP_AM			8'h88
`define OP_AMD			8'h89
`define OP_NM			8'h8a
`define OP_OM			8'h8b
`define OP_XM			8'h8c
`define OP_CM			8'h8d
`define OP_ADC			8'h8e
`define OP_BR7			8'h8f
`define OP_BF			8'h9x
`define OP_INS			8'hax
`define OP_OUTS			8'hbx
`define OP_AS			8'hcx
`define OP_ASD			8'hdx
`define OP_XS			8'hex
`define OP_NS			8'hfx

`define ALU_L		4'h0
`define ALU_R		4'h1
`define ALU_SL_1	4'h2 
`define ALU_SR_1	4'h3
`define ALU_SL_4	4'h4
`define ALU_SR_4	4'h5
`define ALU_LINK	4'h6
`define ALU_COM		4'h7 
`define ALU_INC		4'h8
`define ALU_AND		4'h9
`define ALU_OR		4'ha
`define ALU_XOR		4'hb
`define ALU_ADD		4'hc
`define ALU_CMP		4'hd
`define ALU_ADD_BCD		4'he
`define ALU_DEC_R	4'hf

`endif